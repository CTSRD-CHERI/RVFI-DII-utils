/*-
 * Copyright (c) 2018 Jonathan Woodruff
 * Copyright (c) 2018 Alexandre Joannou
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory (Department of Computer Science and
 * Technology) under DARPA contract HR0011-18-C-0016 ("ECATS"), as part of the
 * DARPA SSITH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 */

import FIFO::*;
import GetPut::*;
import ClientServer::*;
import Connectable :: *;
import RVFI_DII::*;
import RVFI_DII_Bridge::*;

module mkDUT (RVFI_DII_Server);
  FIFO#(RVFI_DII_Execution#(32, 4)) tracebuf <- mkFIFO;
  Reg#(Bit#(64)) count <- mkReg(0);
  interface Put request;
    method put(inst) = action
      tracebuf.enq(RVFI_DII_Execution{
        rvfi_order: count,
        rvfi_trap:  ?,
        rvfi_halt:  ?,
        rvfi_intr:  ?,
        rvfi_insn: inst,
        rvfi_rs1_addr:  ?,
        rvfi_rs2_addr:  ?,
        rvfi_rs1_data:  ?,
        rvfi_rs2_data:  ?,
        rvfi_pc_rdata:  ?,
        rvfi_pc_wdata:  ?,
        rvfi_mem_wdata: ?,
        rvfi_rd_addr:   ?,
        rvfi_rd_wdata:  ?,
        rvfi_mem_addr:  ?,
        rvfi_mem_rmask: ?,
        rvfi_mem_wmask: ?,
        rvfi_mem_rdata: ?
      });
      count <= count + 1;
    endaction;
  endinterface
  interface response = toGet(tracebuf);
endmodule

module mkRVFI_DII_Test(Empty);
  RVFI_DII_Bridge bridge <- mkRVFI_DII_Bridge("RVFI_DII", 5000);
  RVFI_DII_Server    dut <- mkDUT(reset_by bridge.new_rst);
  mkConnection(bridge.inst, dut);
endmodule
